-- Your Names:  Linqiao (James) Liu; Henry Hao Yan
-- Your Student Numbers: 39140116; 59057159
-- Your Lab Section:  L1B

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;